module UpDown(clk, reset, en, s, o);
	parameter n = 4;
	input clk, reset, en, s;
	output reg [n-1:0]o;
	reg initVal = 4'b1010;
	
	initial
		begin
			o = initVal;
		end
		
	always @ (posedge clk)
		begin
			if(!reset)
				begin
					o = initVal;
				end
			else
				begin
					if(!en)
						begin
							o = {n{1'b0}};
						end
					else
						begin
							if(s==0)
								begin
									o = o+1;
								end
							else
								begin
									o = o-1;
								end
						end
				end	
		end
endmodule
