// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 9.1 Build 222 10/21/2009 SJ Full Version
// Created on Tue Apr 16 16:04:09 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module TFF_SD (
    reset,clock,t,
    q);

    input reset;
    input clock;
    input t;
    tri0 reset;
    tri0 t;
    output q;
    reg q;
    reg reg_q;
    reg [1:0] fstate;
    reg [1:0] reg_fstate;
    parameter s0=0,s1=1;

    initial
    begin
        reg_q <= 1'b0;
    end

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or t or reg_q)
    begin
        if (reset) begin
            reg_fstate <= s0;
            reg_q <= 1'b0;
            q <= 1'b0;
        end
        else begin
            reg_q <= 1'b0;
            q <= 1'b0;
            case (fstate)
                s0: begin
                    if (~(t))
                        reg_fstate <= s0;
                    else if (t)
                        reg_fstate <= s1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s0;

                    reg_q <= 1'b0;
                end
                s1: begin
                    if (~(t))
                        reg_fstate <= s1;
                    else if (t)
                        reg_fstate <= s0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= s1;

                    reg_q <= 1'b1;
                end
                default: begin
                    reg_q <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
            q <= reg_q;
        end
    end
endmodule // TFF_SD
